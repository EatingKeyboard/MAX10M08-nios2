
module nios (
	clk_clk,
	reset_reset_n,
	uart_0_rxd,
	uart_0_txd);	

	input		clk_clk;
	input		reset_reset_n;
	input		uart_0_rxd;
	output		uart_0_txd;
endmodule
